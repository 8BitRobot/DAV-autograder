`timescale 1ns/1ns // uncomment this line when you push to the autograder!

module miniALU (
    // TODO: define your input and output ports
    // IMPORTANT: for the autograder to run correctly, you must use the port names we provide
    op1,
    op2, 
    operation,
    sign, 
    result
    );

    // The following block will contain the logic of your combinational circuit
    always_comb begin
        // TODO: write the logic for your miniALU here
    end
endmodule